module mux3 #(parameter WIDTH = 32) (
    input  logic [WIDTH-1:0] a, b, c,
    input  logic [1:0]       sel,
    output logic [WIDTH-1:0] out
);
    always_comb begin
        case (sel)
            2'b00: out = a;
            2'b01: out = b;
            2'b10: out = c;
            default: out = {WIDTH{1'b0}};  // Zero-pad for safety
        endcase
    end
endmodule
